// Type-Parameterized Interface
// testbench
`include "interface.sv"
`include "test.sv"

module testbench;
  intf #(longint, byte) intff();	// initialize  parameter interface
  test tst(intff);		// passing arguments test (test handle)
  
  // instantation with interface to dut
  square dut(intff);
  
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars;
  end
  
endmodule