// Type-Parameterized Interface
// design
module square(intf intff);
  
  assign intff.z = (intff.a ** 2);			// square
endmodule
