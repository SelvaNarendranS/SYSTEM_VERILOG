// interface - simple interface
// interface
interface intf;
  logic a, b;
  logic z;
endinterface